module test;
 wire a,b;
 not A(a,b);
endmodule

