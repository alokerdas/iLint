module test;
`define  WIDTH 128 //warning here
`define  SIZE WIDTH*2 //warning here
`define AA bb
endmodule

