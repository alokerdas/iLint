module TEST; //warning on "TEST_TOP", using
         //"TOP_module" like
endmodule

