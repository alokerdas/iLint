macromodule test( carry, sum, cin, a, b); //non-synthesizable, warning
input carry, a, b;
output sum;
inout cin;
endmodule

