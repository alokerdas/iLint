module test;
 function integer TF; //warning
   input a, b, cin;
   TF = a + b + cin;
 endfunction
endmodule

