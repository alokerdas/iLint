module test;
reg [7:0] mem [0:1023];
endmodule

