module test (A,B,Q,LINE);
input A;
input B; //group input port together
output Q; //separate the ports with different direction by a?
//blank line if the first argument is TRUE.
inout LINE;
endmodule

