module test;
 task Check_0123456789012; //warning on "Check_0123456789012"
 begin
 end
 endtask
endmodule

