module test;
specify
//non-synthesizable, warning here
endspecify
endmodule

