module test;
wire bind,b,c;
and AA(bind,b,c);
endmodule

