module test (a, b, c, d, f);
input a, b, c, d;
output f;
and and1(f, a, b);
or or1(f, c, d);
endmodule

