
module test();
reg signal;
parameter y = 4; 
endmodule

