module test;
 task Check; //warning on "Check"
 begin
 end
 endtask
endmodule

