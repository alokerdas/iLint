`define bytesize 1
`define var_nand(dly) nand #dly
`define wordsize 8
module test (A);
input A;
endmodule
