module test(clock, reset, clock1, reset1, count);
input clock; input reset; //warning here
input clock1;  output reset1;
output count;
endmodule

