module test;
 parameter par_012345678901234 = 5;
       //warning on "par_012345678901234"
endmodule

