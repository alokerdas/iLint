module test(a, b);
 input b;
 output a;
 real c;
 assign a = c;
endmodule

