module test(clock, set, reset, count);
input clock, set;
input reset; //comment
output count;
endmodule
