module test(a,b);
input a;
output b;
not N(b,a);
endmodule

