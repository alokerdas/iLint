//module begin *****OK*******
/*Module
******warning here********
**sub
*/
module sub(clk, i, o);/*sub module*/ //*******warning here*******
input clk, i;
output o;
endmodule

