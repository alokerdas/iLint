module test (a, b, c);
 input a, b;
 output c;
 and and1(c, a, b); //warning on 'and1'
endmodule

