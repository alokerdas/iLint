module test;
wire in,b,c;
and AA(in,b,c);
endmodule

