module test;
 function Func_add;
       //warning on "Func_add"
 input a;
 input b;
 begin
 end
 endfunction
endmodule

