module test;
wire wor_o,b,c;
and AA(wor_o,b,c);
endmodule

