module test;
 function add; //warning on "add", using "f_add" like
 input a;
 input b;
 begin
 end
 endfunction
endmodule

