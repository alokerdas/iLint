module test;
wire export, b, c;
and AA(export, b, c);
endmodule

