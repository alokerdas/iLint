module test;
 task Check; //warning on "Check", using "p_Check" like
 begin
 end
 endtask
endmodule

