module test;
endmodule

