module test(o,a,b,c);
input [8:1]b;
output [9:0]c;
input [0:2] a;
output [3:0] o;
assign o=a;
assign b = c;
endmodule

