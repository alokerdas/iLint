module test;
parameter NOT_OK = 0; // nLint gives warning on this declaration
localparam OK = 1;
endmodule

