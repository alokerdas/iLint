module test(a);
 input a;
 wire a;
 reg b;
endmodule

