module test (clk, d, q, );               
input clk, d;
output q;
//a null port after "q" is used
endmodule
