module test_top_0123456789012;
//warning on "test_top_0123456789012"
endmodule

