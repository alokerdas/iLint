module test1 (o, a);
input a;
output o;
wire b, c;
assign o = c;
assign b = a;
endmodule
