module test;
realtime rt;//non-synthesizable, warning
endmodule

