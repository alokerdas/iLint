module test (A,B,Q,LINE);
input A;
input B; 
output Q; 
inout LINE;
endmodule

