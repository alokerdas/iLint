module TEST_TOP; //warning on "TEST_TOP"
endmodule

