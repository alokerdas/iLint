module test (bind, b, c); //no output for module test
 input bind, b, c;
 and an(bind,b,c);
endmodule

