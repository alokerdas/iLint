module test (clock, q_nxt, q);
 input clock, q_nxt;
 output q;
 reg q;
 always @(posedge clock)
 if(clock)
 begin
 end
endmodule

