module test;
 parameter TW= 33'b100010000000000000000000000000010; //warning here
endmodule

