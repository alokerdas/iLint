module test;
 function real testfun; //warning
   input a, b, cin;
  testfun = a + b + cin;
 endfunction
endmodule

