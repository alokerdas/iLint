module document();
endmodule

