module test;
 wire c;
 reg a,b,d;
 initial
 begin
 assign a=b;
 assign d=c;
 end
endmodule

