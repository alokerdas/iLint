module test (a1234567890123456, b, C);
 input a1234567890123456, b;
 output C;
 wire C;
 and and1(C,a1234567890123456,b);
endmodule

